-- stateMachine_CP_tb